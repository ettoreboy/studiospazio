<?xml version="1.0" encoding="UTF-8"?>
<Batch version="2.0"><TaskList><Task type="OptimizeForWebTask" enabled="True"><FilePath><![CDATA[<Source Folder>]]></FilePath><FileExists>0</FileExists><FileFormat>0</FileFormat><Profile>0</Profile><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGChromaSubsampling>1</JPEGChromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><JPEGRemoveMarkers>False</JPEGRemoveMarkers><JPEGProgressive>True</JPEGProgressive><JPEGBlur>0</JPEGBlur><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGTransparency>True</PNGTransparency><PNGUsePalette>False</PNGUsePalette><PNGColorCount>256</PNGColorCount><PNGInterlaced>False</PNGInterlaced><PNGRemoveTextFields>False</PNGRemoveTextFields><PNGQuality>100</PNGQuality><GIFColorCount>256</GIFColorCount><GIFTransparency>0</GIFTransparency><GIFInterlaced>0</GIFInterlaced><RemoveAllMetadata>0</RemoveAllMetadata></Task></TaskList></Batch>
