<?xml version="1.0" encoding="UTF-8"?>
<Batch version="2.0"><TaskList><Task type="ResizeTask" enabled="True"><Width units="0">-1</Width><Height units="0">1200</Height><DPI>-1</DPI><Filter>8</Filter><UseProportions>True</UseProportions><ResizeType>1</ResizeType></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[1200_<Original Name (Without Extension)>]]></FileName><PreserveStruct>False</PreserveStruct><CommonFolder><![CDATA[]]></CommonFolder><FileType></FileType><FilePath><![CDATA[<Source Folder>]]></FilePath><FileExists>1</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed><DDSMIPLevels>8</DDSMIPLevels><DDSMipMapFilter>4</DDSMipMapFilter><DDSFormat>71</DDSFormat></Task><Task type="ResizeTask" enabled="True"><Width units="0">-1</Width><Height units="0">768</Height><DPI>-1</DPI><Filter>8</Filter><UseProportions>True</UseProportions><ResizeType>1</ResizeType></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[768_<Original Name (Without Extension)>]]></FileName><PreserveStruct>False</PreserveStruct><CommonFolder><![CDATA[]]></CommonFolder><FileType>JPEG</FileType><FilePath><![CDATA[<Source Folder>]]></FilePath><FileExists>1</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed><DDSMIPLevels>8</DDSMIPLevels><DDSMipMapFilter>4</DDSMipMapFilter><DDSFormat>71</DDSFormat></Task><Task type="ResizeTask" enabled="True"><Width units="0">480</Width><Height units="0">-1</Height><DPI>-1</DPI><Filter>8</Filter><UseProportions>True</UseProportions><ResizeType>1</ResizeType></Task></TaskList></Batch>
