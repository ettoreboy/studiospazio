<?xml version="1.0" encoding="UTF-8"?>
<Batch version="2.0"><TaskList><Task type="FileCopyTask" enabled="True"><FileName><![CDATA[orig_<Original Name (Without Extension)>]]></FileName><FilePath><![CDATA[<Source Folder>]]></FilePath><PreserveStructure>0</PreserveStructure><CommonFolder><![CDATA[C:\Users\ciprian\Documents\GitHub\studiospazio\projects\1_GarageSuzzara\]]></CommonFolder><FileExists>3</FileExists></Task><Task type="ResizeTask" enabled="True"><Width units="0">-1</Width><Height units="0">1050</Height><DPI>-1</DPI><Filter>8</Filter><UseProportions>True</UseProportions><ResizeType>0</ResizeType></Task><Task type="FileCopyTask" enabled="True"><FileName><![CDATA[1050_<Original Name (Without Extension)>]]></FileName><FilePath><![CDATA[<Source Folder>]]></FilePath><PreserveStructure>0</PreserveStructure><CommonFolder><![CDATA[C:\Users\ciprian\Documents\GitHub\studiospazio\projects\1_GarageSuzzara\]]></CommonFolder><FileExists>0</FileExists></Task><Task type="ResizeTask" enabled="True"><Width units="0">-1</Width><Height units="0">720</Height><DPI>-1</DPI><Filter>8</Filter><UseProportions>True</UseProportions><ResizeType>0</ResizeType></Task><Task type="FileCopyTask" enabled="True"><FileName><![CDATA[720_<Original Name (Without Extension)>]]></FileName><FilePath><![CDATA[<Source Folder>]]></FilePath><PreserveStructure>0</PreserveStructure><CommonFolder><![CDATA[C:\Users\ciprian\Documents\GitHub\studiospazio\projects\1_GarageSuzzara\]]></CommonFolder><FileExists>0</FileExists></Task><Task type="ResizeTask" enabled="True"><Width units="0">480</Width><Height units="0">-1</Height><DPI>-1</DPI><Filter>8</Filter><UseProportions>True</UseProportions><ResizeType>0</ResizeType></Task><Task type="RenameTask" enabled="True"><FileName><![CDATA[480_<Original Name (Without Extension)>]]></FileName><FilePath><![CDATA[<Source Folder>]]></FilePath><PreserveStruct>0</PreserveStruct><CommonFolder><![CDATA[]]></CommonFolder><FileExists>3</FileExists><Cases>0</Cases></Task><Task type="OptimizeForWebTask" enabled="True"><FilePath><![CDATA[<Source Folder>]]></FilePath><FileExists>3</FileExists><FileFormat>0</FileFormat><Profile>0</Profile><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGChromaSubsampling>1</JPEGChromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><JPEGRemoveMarkers>False</JPEGRemoveMarkers><JPEGProgressive>False</JPEGProgressive><JPEGBlur>0</JPEGBlur><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGTransparency>True</PNGTransparency><PNGUsePalette>False</PNGUsePalette><PNGColorCount>256</PNGColorCount><PNGInterlaced>False</PNGInterlaced><PNGRemoveTextFields>False</PNGRemoveTextFields><PNGQuality>100</PNGQuality><GIFColorCount>256</GIFColorCount><GIFTransparency>0</GIFTransparency><GIFInterlaced>0</GIFInterlaced><RemoveAllMetadata>0</RemoveAllMetadata></Task></TaskList></Batch>
